// nios.v

// Generated using ACDS version 17.0 602

`timescale 1 ps / 1 ps
module nios (
		input  wire       busy_export,     //     busy.export
		output wire [9:0] bx_export,       //       bx.export
		output wire [9:0] by_export,       //       by.export
		input  wire       clk_clk,         //      clk.clk
		output wire       lcd_out_rs,      //  lcd_out.rs
		output wire       lcd_out_rw,      //         .rw
		output wire       lcd_out_en,      //         .en
		output wire [7:0] lcd_out_db,      //         .db
		output wire [9:0] p1x_export,      //      p1x.export
		output wire [9:0] p1y_export,      //      p1y.export
		output wire [9:0] p2x_export,      //      p2x.export
		output wire [9:0] p2y_export,      //      p2y.export
		input  wire [7:0] player1_export,  //  player1.export
		input  wire [7:0] player_2_export, // player_2.export
		input  wire       reset_reset_n,   //    reset.reset_n
		input  wire       start_export     //    start.export
	);

	wire         nios_custom_instruction_master_readra;                                   // nios:D_ci_readra -> nios_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_a;                                        // nios:D_ci_a -> nios_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_b;                                        // nios:D_ci_b -> nios_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_c;                                        // nios:D_ci_c -> nios_custom_instruction_master_translator:ci_slave_c
	wire         nios_custom_instruction_master_readrb;                                   // nios:D_ci_readrb -> nios_custom_instruction_master_translator:ci_slave_readrb
	wire         nios_custom_instruction_master_clk;                                      // nios:E_ci_multi_clock -> nios_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios_custom_instruction_master_ipending;                                 // nios:W_ci_ipending -> nios_custom_instruction_master_translator:ci_slave_ipending
	wire         nios_custom_instruction_master_start;                                    // nios:E_ci_multi_start -> nios_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios_custom_instruction_master_reset_req;                                // nios:E_ci_multi_reset_req -> nios_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios_custom_instruction_master_done;                                     // nios_custom_instruction_master_translator:ci_slave_multi_done -> nios:E_ci_multi_done
	wire   [7:0] nios_custom_instruction_master_n;                                        // nios:D_ci_n -> nios_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_result;                                   // nios_custom_instruction_master_translator:ci_slave_result -> nios:E_ci_result
	wire         nios_custom_instruction_master_estatus;                                  // nios:W_ci_estatus -> nios_custom_instruction_master_translator:ci_slave_estatus
	wire         nios_custom_instruction_master_clk_en;                                   // nios:E_ci_multi_clk_en -> nios_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] nios_custom_instruction_master_datab;                                    // nios:E_ci_datab -> nios_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_dataa;                                    // nios:E_ci_dataa -> nios_custom_instruction_master_translator:ci_slave_dataa
	wire         nios_custom_instruction_master_reset;                                    // nios:E_ci_multi_reset -> nios_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios_custom_instruction_master_writerc;                                  // nios:D_ci_writerc -> nios_custom_instruction_master_translator:ci_slave_writerc
	wire         nios_custom_instruction_master_translator_multi_ci_master_readra;        // nios_custom_instruction_master_translator:multi_ci_master_readra -> nios_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_a;             // nios_custom_instruction_master_translator:multi_ci_master_a -> nios_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_b;             // nios_custom_instruction_master_translator:multi_ci_master_b -> nios_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk;           // nios_custom_instruction_master_translator:multi_ci_master_clk -> nios_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios_custom_instruction_master_translator_multi_ci_master_readrb;        // nios_custom_instruction_master_translator:multi_ci_master_readrb -> nios_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_c;             // nios_custom_instruction_master_translator:multi_ci_master_c -> nios_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios_custom_instruction_master_translator_multi_ci_master_start;         // nios_custom_instruction_master_translator:multi_ci_master_start -> nios_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios_custom_instruction_master_translator:multi_ci_master_reset_req -> nios_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios_custom_instruction_master_translator_multi_ci_master_done;          // nios_custom_instruction_master_multi_xconnect:ci_slave_done -> nios_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios_custom_instruction_master_translator_multi_ci_master_n;             // nios_custom_instruction_master_translator:multi_ci_master_n -> nios_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_result;        // nios_custom_instruction_master_multi_xconnect:ci_slave_result -> nios_custom_instruction_master_translator:multi_ci_master_result
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios_custom_instruction_master_translator:multi_ci_master_clken -> nios_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_datab;         // nios_custom_instruction_master_translator:multi_ci_master_datab -> nios_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_dataa;         // nios_custom_instruction_master_translator:multi_ci_master_dataa -> nios_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset;         // nios_custom_instruction_master_translator:multi_ci_master_reset -> nios_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios_custom_instruction_master_translator_multi_ci_master_writerc;       // nios_custom_instruction_master_translator:multi_ci_master_writerc -> nios_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios_custom_instruction_master_multi_xconnect:ci_master0_a -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios_custom_instruction_master_multi_xconnect:ci_master0_b -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios_custom_instruction_master_multi_xconnect:ci_master0_c -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios_custom_instruction_master_multi_xconnect:ci_master0_start -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios_custom_instruction_master_multi_xconnect:ci_master0_n -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_result; // delay_0:result -> nios_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios_custom_instruction_master_multi_slave_translator0:ci_master_clk -> delay_0:clk
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios_custom_instruction_master_multi_slave_translator0:ci_master_clken -> delay_0:clk_en
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_datab -> delay_0:datab
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> delay_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_start -> delay_0:start
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_reset -> delay_0:reset
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_done;   // delay_0:done -> nios_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios_custom_instruction_master_multi_xconnect:ci_master1_a -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios_custom_instruction_master_multi_xconnect:ci_master1_b -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios_custom_instruction_master_multi_xconnect:ci_master1_c -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios_custom_instruction_master_multi_xconnect:ci_master1_start -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios_custom_instruction_master_multi_xconnect:ci_master1_n -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator1_ci_master_result; // div_0:result -> nios_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios_custom_instruction_master_multi_slave_translator1:ci_master_clk -> div_0:clk
	wire         nios_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios_custom_instruction_master_multi_slave_translator1:ci_master_clken -> div_0:clk_en
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // nios_custom_instruction_master_multi_slave_translator1:ci_master_datab -> div_0:datab
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> div_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator1_ci_master_start;  // nios_custom_instruction_master_multi_slave_translator1:ci_master_start -> div_0:start
	wire         nios_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios_custom_instruction_master_multi_slave_translator1:ci_master_reset -> div_0:reset
	wire         nios_custom_instruction_master_multi_slave_translator1_ci_master_done;   // div_0:done -> nios_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_readra;         // nios_custom_instruction_master_multi_xconnect:ci_master2_readra -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master2_a;              // nios_custom_instruction_master_multi_xconnect:ci_master2_a -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master2_b;              // nios_custom_instruction_master_multi_xconnect:ci_master2_b -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_b
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_readrb;         // nios_custom_instruction_master_multi_xconnect:ci_master2_readrb -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_readrb
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master2_c;              // nios_custom_instruction_master_multi_xconnect:ci_master2_c -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_clk;            // nios_custom_instruction_master_multi_xconnect:ci_master2_clk -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_clk
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master2_ipending;       // nios_custom_instruction_master_multi_xconnect:ci_master2_ipending -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_start;          // nios_custom_instruction_master_multi_xconnect:ci_master2_start -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_start
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_reset_req;      // nios_custom_instruction_master_multi_xconnect:ci_master2_reset_req -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_done;           // nios_custom_instruction_master_multi_slave_translator2:ci_slave_done -> nios_custom_instruction_master_multi_xconnect:ci_master2_done
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master2_n;              // nios_custom_instruction_master_multi_xconnect:ci_master2_n -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master2_result;         // nios_custom_instruction_master_multi_slave_translator2:ci_slave_result -> nios_custom_instruction_master_multi_xconnect:ci_master2_result
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_estatus;        // nios_custom_instruction_master_multi_xconnect:ci_master2_estatus -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_estatus
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_clk_en;         // nios_custom_instruction_master_multi_xconnect:ci_master2_clken -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_clken
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master2_datab;          // nios_custom_instruction_master_multi_xconnect:ci_master2_datab -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master2_dataa;          // nios_custom_instruction_master_multi_xconnect:ci_master2_dataa -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_reset;          // nios_custom_instruction_master_multi_xconnect:ci_master2_reset -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_reset
	wire         nios_custom_instruction_master_multi_xconnect_ci_master2_writerc;        // nios_custom_instruction_master_multi_xconnect:ci_master2_writerc -> nios_custom_instruction_master_multi_slave_translator2:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator2_ci_master_result; // lcd_0:result -> nios_custom_instruction_master_multi_slave_translator2:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator2_ci_master_clk;    // nios_custom_instruction_master_multi_slave_translator2:ci_master_clk -> lcd_0:clk
	wire         nios_custom_instruction_master_multi_slave_translator2_ci_master_clk_en; // nios_custom_instruction_master_multi_slave_translator2:ci_master_clken -> lcd_0:clk_en
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator2_ci_master_datab;  // nios_custom_instruction_master_multi_slave_translator2:ci_master_datab -> lcd_0:datab
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator2_ci_master_dataa;  // nios_custom_instruction_master_multi_slave_translator2:ci_master_dataa -> lcd_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator2_ci_master_start;  // nios_custom_instruction_master_multi_slave_translator2:ci_master_start -> lcd_0:start
	wire         nios_custom_instruction_master_multi_slave_translator2_ci_master_reset;  // nios_custom_instruction_master_multi_slave_translator2:ci_master_reset -> lcd_0:reset
	wire         nios_custom_instruction_master_multi_slave_translator2_ci_master_done;   // lcd_0:done -> nios_custom_instruction_master_multi_slave_translator2:ci_master_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_readra;         // nios_custom_instruction_master_multi_xconnect:ci_master3_readra -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_readra
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master3_a;              // nios_custom_instruction_master_multi_xconnect:ci_master3_a -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_a
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master3_b;              // nios_custom_instruction_master_multi_xconnect:ci_master3_b -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_b
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_readrb;         // nios_custom_instruction_master_multi_xconnect:ci_master3_readrb -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_readrb
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master3_c;              // nios_custom_instruction_master_multi_xconnect:ci_master3_c -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_clk;            // nios_custom_instruction_master_multi_xconnect:ci_master3_clk -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_clk
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master3_ipending;       // nios_custom_instruction_master_multi_xconnect:ci_master3_ipending -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_start;          // nios_custom_instruction_master_multi_xconnect:ci_master3_start -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_start
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_reset_req;      // nios_custom_instruction_master_multi_xconnect:ci_master3_reset_req -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_done;           // nios_custom_instruction_master_multi_slave_translator3:ci_slave_done -> nios_custom_instruction_master_multi_xconnect:ci_master3_done
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master3_n;              // nios_custom_instruction_master_multi_xconnect:ci_master3_n -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_n
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master3_result;         // nios_custom_instruction_master_multi_slave_translator3:ci_slave_result -> nios_custom_instruction_master_multi_xconnect:ci_master3_result
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_estatus;        // nios_custom_instruction_master_multi_xconnect:ci_master3_estatus -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_estatus
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_clk_en;         // nios_custom_instruction_master_multi_xconnect:ci_master3_clken -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_clken
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master3_datab;          // nios_custom_instruction_master_multi_xconnect:ci_master3_datab -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_datab
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master3_dataa;          // nios_custom_instruction_master_multi_xconnect:ci_master3_dataa -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_reset;          // nios_custom_instruction_master_multi_xconnect:ci_master3_reset -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_reset
	wire         nios_custom_instruction_master_multi_xconnect_ci_master3_writerc;        // nios_custom_instruction_master_multi_xconnect:ci_master3_writerc -> nios_custom_instruction_master_multi_slave_translator3:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator3_ci_master_result; // mult:result -> nios_custom_instruction_master_multi_slave_translator3:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator3_ci_master_clk;    // nios_custom_instruction_master_multi_slave_translator3:ci_master_clk -> mult:clk
	wire         nios_custom_instruction_master_multi_slave_translator3_ci_master_clk_en; // nios_custom_instruction_master_multi_slave_translator3:ci_master_clken -> mult:clk_en
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator3_ci_master_datab;  // nios_custom_instruction_master_multi_slave_translator3:ci_master_datab -> mult:datab
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator3_ci_master_dataa;  // nios_custom_instruction_master_multi_slave_translator3:ci_master_dataa -> mult:dataa
	wire         nios_custom_instruction_master_multi_slave_translator3_ci_master_start;  // nios_custom_instruction_master_multi_slave_translator3:ci_master_start -> mult:start
	wire         nios_custom_instruction_master_multi_slave_translator3_ci_master_reset;  // nios_custom_instruction_master_multi_slave_translator3:ci_master_reset -> mult:reset
	wire         nios_custom_instruction_master_multi_slave_translator3_ci_master_done;   // mult:done -> nios_custom_instruction_master_multi_slave_translator3:ci_master_done
	wire  [31:0] nios_data_master_readdata;                                               // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                                            // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                                            // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [14:0] nios_data_master_address;                                                // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                                             // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                                   // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                                                  // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                              // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                                        // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                                     // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [14:0] nios_instruction_master_address;                                         // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                                            // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;                         // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;                      // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;                          // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;                             // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;                            // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;                        // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                                  // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                    // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire  [10:0] mm_interconnect_0_memory_s1_address;                                     // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                  // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                                       // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                   // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                                       // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire  [31:0] mm_interconnect_0_start_s1_readdata;                                     // start:readdata -> mm_interconnect_0:start_s1_readdata
	wire   [1:0] mm_interconnect_0_start_s1_address;                                      // mm_interconnect_0:start_s1_address -> start:address
	wire         mm_interconnect_0_p1x_s1_chipselect;                                     // mm_interconnect_0:p1x_s1_chipselect -> p1x:chipselect
	wire  [31:0] mm_interconnect_0_p1x_s1_readdata;                                       // p1x:readdata -> mm_interconnect_0:p1x_s1_readdata
	wire   [1:0] mm_interconnect_0_p1x_s1_address;                                        // mm_interconnect_0:p1x_s1_address -> p1x:address
	wire         mm_interconnect_0_p1x_s1_write;                                          // mm_interconnect_0:p1x_s1_write -> p1x:write_n
	wire  [31:0] mm_interconnect_0_p1x_s1_writedata;                                      // mm_interconnect_0:p1x_s1_writedata -> p1x:writedata
	wire         mm_interconnect_0_p1y_s1_chipselect;                                     // mm_interconnect_0:p1y_s1_chipselect -> p1y:chipselect
	wire  [31:0] mm_interconnect_0_p1y_s1_readdata;                                       // p1y:readdata -> mm_interconnect_0:p1y_s1_readdata
	wire   [1:0] mm_interconnect_0_p1y_s1_address;                                        // mm_interconnect_0:p1y_s1_address -> p1y:address
	wire         mm_interconnect_0_p1y_s1_write;                                          // mm_interconnect_0:p1y_s1_write -> p1y:write_n
	wire  [31:0] mm_interconnect_0_p1y_s1_writedata;                                      // mm_interconnect_0:p1y_s1_writedata -> p1y:writedata
	wire         mm_interconnect_0_p2x_s1_chipselect;                                     // mm_interconnect_0:p2x_s1_chipselect -> p2x:chipselect
	wire  [31:0] mm_interconnect_0_p2x_s1_readdata;                                       // p2x:readdata -> mm_interconnect_0:p2x_s1_readdata
	wire   [1:0] mm_interconnect_0_p2x_s1_address;                                        // mm_interconnect_0:p2x_s1_address -> p2x:address
	wire         mm_interconnect_0_p2x_s1_write;                                          // mm_interconnect_0:p2x_s1_write -> p2x:write_n
	wire  [31:0] mm_interconnect_0_p2x_s1_writedata;                                      // mm_interconnect_0:p2x_s1_writedata -> p2x:writedata
	wire         mm_interconnect_0_p2y_s1_chipselect;                                     // mm_interconnect_0:p2y_s1_chipselect -> p2y:chipselect
	wire  [31:0] mm_interconnect_0_p2y_s1_readdata;                                       // p2y:readdata -> mm_interconnect_0:p2y_s1_readdata
	wire   [1:0] mm_interconnect_0_p2y_s1_address;                                        // mm_interconnect_0:p2y_s1_address -> p2y:address
	wire         mm_interconnect_0_p2y_s1_write;                                          // mm_interconnect_0:p2y_s1_write -> p2y:write_n
	wire  [31:0] mm_interconnect_0_p2y_s1_writedata;                                      // mm_interconnect_0:p2y_s1_writedata -> p2y:writedata
	wire         mm_interconnect_0_bx_s1_chipselect;                                      // mm_interconnect_0:bx_s1_chipselect -> bx:chipselect
	wire  [31:0] mm_interconnect_0_bx_s1_readdata;                                        // bx:readdata -> mm_interconnect_0:bx_s1_readdata
	wire   [1:0] mm_interconnect_0_bx_s1_address;                                         // mm_interconnect_0:bx_s1_address -> bx:address
	wire         mm_interconnect_0_bx_s1_write;                                           // mm_interconnect_0:bx_s1_write -> bx:write_n
	wire  [31:0] mm_interconnect_0_bx_s1_writedata;                                       // mm_interconnect_0:bx_s1_writedata -> bx:writedata
	wire         mm_interconnect_0_by_s1_chipselect;                                      // mm_interconnect_0:by_s1_chipselect -> by:chipselect
	wire  [31:0] mm_interconnect_0_by_s1_readdata;                                        // by:readdata -> mm_interconnect_0:by_s1_readdata
	wire   [1:0] mm_interconnect_0_by_s1_address;                                         // mm_interconnect_0:by_s1_address -> by:address
	wire         mm_interconnect_0_by_s1_write;                                           // mm_interconnect_0:by_s1_write -> by:write_n
	wire  [31:0] mm_interconnect_0_by_s1_writedata;                                       // mm_interconnect_0:by_s1_writedata -> by:writedata
	wire  [31:0] mm_interconnect_0_player1_s1_readdata;                                   // player1:readdata -> mm_interconnect_0:player1_s1_readdata
	wire   [1:0] mm_interconnect_0_player1_s1_address;                                    // mm_interconnect_0:player1_s1_address -> player1:address
	wire  [31:0] mm_interconnect_0_player_2_s1_readdata;                                  // player_2:readdata -> mm_interconnect_0:player_2_s1_readdata
	wire   [1:0] mm_interconnect_0_player_2_s1_address;                                   // mm_interconnect_0:player_2_s1_address -> player_2:address
	wire  [31:0] mm_interconnect_0_busy_s1_readdata;                                      // busy:readdata -> mm_interconnect_0:busy_s1_readdata
	wire   [1:0] mm_interconnect_0_busy_s1_address;                                       // mm_interconnect_0:busy_s1_address -> busy:address
	wire  [31:0] nios_irq_irq;                                                            // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [busy:reset_n, bx:reset_n, by:reset_n, irq_mapper:reset, memory:reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, p1x:reset_n, p1y:reset_n, p2x:reset_n, p2y:reset_n, player1:reset_n, player_2:reset_n, rst_translator:in_reset, start:reset_n]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [memory:reset_req, nios:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                                          // nios:debug_reset_request -> rst_controller:reset_in1

	nios_busy busy (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_busy_s1_readdata), //                    .readdata
		.in_port  (busy_export)                         // external_connection.export
	);

	nios_bx bx (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_bx_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bx_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bx_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bx_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bx_s1_readdata),   //                    .readdata
		.out_port   (bx_export)                           // external_connection.export
	);

	nios_bx by (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_by_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_by_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_by_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_by_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_by_s1_readdata),   //                    .readdata
		.out_port   (by_export)                           // external_connection.export
	);

	delay30fps delay_0 (
		.dataa  (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // delay_instr.dataa
		.datab  (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //            .datab
		.result (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //            .result
		.clk    (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //            .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //            .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //            .start
		.reset  (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //            .reset
		.done   (nios_custom_instruction_master_multi_slave_translator0_ci_master_done)    //            .done
	);

	div div_0 (
		.reset  (nios_custom_instruction_master_multi_slave_translator1_ci_master_reset),  // div_instr.reset
		.clk    (nios_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.done   (nios_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.start  (nios_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.clk_en (nios_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.result (nios_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.datab  (nios_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.dataa  (nios_custom_instruction_master_multi_slave_translator1_ci_master_dataa)   //          .dataa
	);

	lcd_driver lcd_0 (
		.dataa  (nios_custom_instruction_master_multi_slave_translator2_ci_master_dataa),  //   lcd_instr.dataa
		.datab  (nios_custom_instruction_master_multi_slave_translator2_ci_master_datab),  //            .datab
		.result (nios_custom_instruction_master_multi_slave_translator2_ci_master_result), //            .result
		.clk    (nios_custom_instruction_master_multi_slave_translator2_ci_master_clk),    //            .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator2_ci_master_clk_en), //            .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator2_ci_master_start),  //            .start
		.reset  (nios_custom_instruction_master_multi_slave_translator2_ci_master_reset),  //            .reset
		.done   (nios_custom_instruction_master_multi_slave_translator2_ci_master_done),   //            .done
		.rs     (lcd_out_rs),                                                              // conduit_lcd.rs
		.rw     (lcd_out_rw),                                                              //            .rw
		.en     (lcd_out_en),                                                              //            .en
		.db     (lcd_out_db)                                                               //            .db
	);

	nios_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	mul mult (
		.dataa  (nios_custom_instruction_master_multi_slave_translator3_ci_master_dataa),  // mult_instr.dataa
		.datab  (nios_custom_instruction_master_multi_slave_translator3_ci_master_datab),  //           .datab
		.result (nios_custom_instruction_master_multi_slave_translator3_ci_master_result), //           .result
		.clk    (nios_custom_instruction_master_multi_slave_translator3_ci_master_clk),    //           .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator3_ci_master_clk_en), //           .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator3_ci_master_start),  //           .start
		.reset  (nios_custom_instruction_master_multi_slave_translator3_ci_master_reset),  //           .reset
		.done   (nios_custom_instruction_master_multi_slave_translator3_ci_master_done)    //           .done
	);

	nios_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (nios_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (nios_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (nios_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (nios_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (nios_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (nios_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (nios_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (nios_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (nios_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios_custom_instruction_master_ipending)             //                          .ipending
	);

	nios_bx p1x (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_p1x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1x_s1_readdata),   //                    .readdata
		.out_port   (p1x_export)                           // external_connection.export
	);

	nios_bx p1y (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_p1y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p1y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p1y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p1y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p1y_s1_readdata),   //                    .readdata
		.out_port   (p1y_export)                           // external_connection.export
	);

	nios_bx p2x (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_p2x_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p2x_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p2x_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p2x_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p2x_s1_readdata),   //                    .readdata
		.out_port   (p2x_export)                           // external_connection.export
	);

	nios_bx p2y (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_p2y_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_p2y_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_p2y_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_p2y_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_p2y_s1_readdata),   //                    .readdata
		.out_port   (p2y_export)                           // external_connection.export
	);

	nios_player1 player1 (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_player1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_player1_s1_readdata), //                    .readdata
		.in_port  (player1_export)                         // external_connection.export
	);

	nios_player1 player_2 (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_player_2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_player_2_s1_readdata), //                    .readdata
		.in_port  (player_2_export)                         // external_connection.export
	);

	nios_busy start (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_start_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_start_s1_readdata), //                    .readdata
		.in_port  (start_export)                         // external_connection.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                    //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                    //                .datab
		.comb_ci_master_result     (),                                                                    //                .result
		.comb_ci_master_n          (),                                                                    //                .n
		.comb_ci_master_readra     (),                                                                    //                .readra
		.comb_ci_master_readrb     (),                                                                    //                .readrb
		.comb_ci_master_writerc    (),                                                                    //                .writerc
		.comb_ci_master_a          (),                                                                    //                .a
		.comb_ci_master_b          (),                                                                    //                .b
		.comb_ci_master_c          (),                                                                    //                .c
		.comb_ci_master_ipending   (),                                                                    //                .ipending
		.comb_ci_master_estatus    (),                                                                    //                .estatus
		.multi_ci_master_clk       (nios_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_result     (),                                                                    //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                         //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                             //     (terminated)
	);

	nios_nios_custom_instruction_master_multi_xconnect nios_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (nios_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios_custom_instruction_master_multi_xconnect_ci_master1_done),       //           .done
		.ci_master2_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master2_dataa),      // ci_master2.dataa
		.ci_master2_datab     (nios_custom_instruction_master_multi_xconnect_ci_master2_datab),      //           .datab
		.ci_master2_result    (nios_custom_instruction_master_multi_xconnect_ci_master2_result),     //           .result
		.ci_master2_n         (nios_custom_instruction_master_multi_xconnect_ci_master2_n),          //           .n
		.ci_master2_readra    (nios_custom_instruction_master_multi_xconnect_ci_master2_readra),     //           .readra
		.ci_master2_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master2_readrb),     //           .readrb
		.ci_master2_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master2_writerc),    //           .writerc
		.ci_master2_a         (nios_custom_instruction_master_multi_xconnect_ci_master2_a),          //           .a
		.ci_master2_b         (nios_custom_instruction_master_multi_xconnect_ci_master2_b),          //           .b
		.ci_master2_c         (nios_custom_instruction_master_multi_xconnect_ci_master2_c),          //           .c
		.ci_master2_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master2_ipending),   //           .ipending
		.ci_master2_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master2_estatus),    //           .estatus
		.ci_master2_clk       (nios_custom_instruction_master_multi_xconnect_ci_master2_clk),        //           .clk
		.ci_master2_reset     (nios_custom_instruction_master_multi_xconnect_ci_master2_reset),      //           .reset
		.ci_master2_clken     (nios_custom_instruction_master_multi_xconnect_ci_master2_clk_en),     //           .clk_en
		.ci_master2_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master2_reset_req),  //           .reset_req
		.ci_master2_start     (nios_custom_instruction_master_multi_xconnect_ci_master2_start),      //           .start
		.ci_master2_done      (nios_custom_instruction_master_multi_xconnect_ci_master2_done),       //           .done
		.ci_master3_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master3_dataa),      // ci_master3.dataa
		.ci_master3_datab     (nios_custom_instruction_master_multi_xconnect_ci_master3_datab),      //           .datab
		.ci_master3_result    (nios_custom_instruction_master_multi_xconnect_ci_master3_result),     //           .result
		.ci_master3_n         (nios_custom_instruction_master_multi_xconnect_ci_master3_n),          //           .n
		.ci_master3_readra    (nios_custom_instruction_master_multi_xconnect_ci_master3_readra),     //           .readra
		.ci_master3_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master3_readrb),     //           .readrb
		.ci_master3_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master3_writerc),    //           .writerc
		.ci_master3_a         (nios_custom_instruction_master_multi_xconnect_ci_master3_a),          //           .a
		.ci_master3_b         (nios_custom_instruction_master_multi_xconnect_ci_master3_b),          //           .b
		.ci_master3_c         (nios_custom_instruction_master_multi_xconnect_ci_master3_c),          //           .c
		.ci_master3_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master3_ipending),   //           .ipending
		.ci_master3_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master3_estatus),    //           .estatus
		.ci_master3_clk       (nios_custom_instruction_master_multi_xconnect_ci_master3_clk),        //           .clk
		.ci_master3_reset     (nios_custom_instruction_master_multi_xconnect_ci_master3_reset),      //           .reset
		.ci_master3_clken     (nios_custom_instruction_master_multi_xconnect_ci_master3_clk_en),     //           .clk_en
		.ci_master3_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master3_reset_req),  //           .reset_req
		.ci_master3_start     (nios_custom_instruction_master_multi_xconnect_ci_master3_start),      //           .start
		.ci_master3_done      (nios_custom_instruction_master_multi_xconnect_ci_master3_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator2 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master2_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master2_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master2_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master2_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master2_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master2_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master2_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master2_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master2_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master2_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master2_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master2_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master2_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master2_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master2_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master2_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master2_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master2_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator2_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator2_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator2_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator2_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator2_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator2_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator2_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator2_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator3 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master3_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master3_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master3_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master3_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master3_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master3_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master3_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master3_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master3_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master3_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master3_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master3_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master3_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master3_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master3_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master3_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master3_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master3_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator3_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator3_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator3_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator3_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator3_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator3_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator3_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator3_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                            (clk_clk),                                            //                          clk_clk.clk
		.nios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address               (nios_data_master_address),                           //                 nios_data_master.address
		.nios_data_master_waitrequest           (nios_data_master_waitrequest),                       //                                 .waitrequest
		.nios_data_master_byteenable            (nios_data_master_byteenable),                        //                                 .byteenable
		.nios_data_master_read                  (nios_data_master_read),                              //                                 .read
		.nios_data_master_readdata              (nios_data_master_readdata),                          //                                 .readdata
		.nios_data_master_write                 (nios_data_master_write),                             //                                 .write
		.nios_data_master_writedata             (nios_data_master_writedata),                         //                                 .writedata
		.nios_data_master_debugaccess           (nios_data_master_debugaccess),                       //                                 .debugaccess
		.nios_instruction_master_address        (nios_instruction_master_address),                    //          nios_instruction_master.address
		.nios_instruction_master_waitrequest    (nios_instruction_master_waitrequest),                //                                 .waitrequest
		.nios_instruction_master_read           (nios_instruction_master_read),                       //                                 .read
		.nios_instruction_master_readdata       (nios_instruction_master_readdata),                   //                                 .readdata
		.busy_s1_address                        (mm_interconnect_0_busy_s1_address),                  //                          busy_s1.address
		.busy_s1_readdata                       (mm_interconnect_0_busy_s1_readdata),                 //                                 .readdata
		.bx_s1_address                          (mm_interconnect_0_bx_s1_address),                    //                            bx_s1.address
		.bx_s1_write                            (mm_interconnect_0_bx_s1_write),                      //                                 .write
		.bx_s1_readdata                         (mm_interconnect_0_bx_s1_readdata),                   //                                 .readdata
		.bx_s1_writedata                        (mm_interconnect_0_bx_s1_writedata),                  //                                 .writedata
		.bx_s1_chipselect                       (mm_interconnect_0_bx_s1_chipselect),                 //                                 .chipselect
		.by_s1_address                          (mm_interconnect_0_by_s1_address),                    //                            by_s1.address
		.by_s1_write                            (mm_interconnect_0_by_s1_write),                      //                                 .write
		.by_s1_readdata                         (mm_interconnect_0_by_s1_readdata),                   //                                 .readdata
		.by_s1_writedata                        (mm_interconnect_0_by_s1_writedata),                  //                                 .writedata
		.by_s1_chipselect                       (mm_interconnect_0_by_s1_chipselect),                 //                                 .chipselect
		.memory_s1_address                      (mm_interconnect_0_memory_s1_address),                //                        memory_s1.address
		.memory_s1_write                        (mm_interconnect_0_memory_s1_write),                  //                                 .write
		.memory_s1_readdata                     (mm_interconnect_0_memory_s1_readdata),               //                                 .readdata
		.memory_s1_writedata                    (mm_interconnect_0_memory_s1_writedata),              //                                 .writedata
		.memory_s1_byteenable                   (mm_interconnect_0_memory_s1_byteenable),             //                                 .byteenable
		.memory_s1_chipselect                   (mm_interconnect_0_memory_s1_chipselect),             //                                 .chipselect
		.memory_s1_clken                        (mm_interconnect_0_memory_s1_clken),                  //                                 .clken
		.nios_debug_mem_slave_address           (mm_interconnect_0_nios_debug_mem_slave_address),     //             nios_debug_mem_slave.address
		.nios_debug_mem_slave_write             (mm_interconnect_0_nios_debug_mem_slave_write),       //                                 .write
		.nios_debug_mem_slave_read              (mm_interconnect_0_nios_debug_mem_slave_read),        //                                 .read
		.nios_debug_mem_slave_readdata          (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                                 .readdata
		.nios_debug_mem_slave_writedata         (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                                 .writedata
		.nios_debug_mem_slave_byteenable        (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                                 .byteenable
		.nios_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                                 .waitrequest
		.nios_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                                 .debugaccess
		.p1x_s1_address                         (mm_interconnect_0_p1x_s1_address),                   //                           p1x_s1.address
		.p1x_s1_write                           (mm_interconnect_0_p1x_s1_write),                     //                                 .write
		.p1x_s1_readdata                        (mm_interconnect_0_p1x_s1_readdata),                  //                                 .readdata
		.p1x_s1_writedata                       (mm_interconnect_0_p1x_s1_writedata),                 //                                 .writedata
		.p1x_s1_chipselect                      (mm_interconnect_0_p1x_s1_chipselect),                //                                 .chipselect
		.p1y_s1_address                         (mm_interconnect_0_p1y_s1_address),                   //                           p1y_s1.address
		.p1y_s1_write                           (mm_interconnect_0_p1y_s1_write),                     //                                 .write
		.p1y_s1_readdata                        (mm_interconnect_0_p1y_s1_readdata),                  //                                 .readdata
		.p1y_s1_writedata                       (mm_interconnect_0_p1y_s1_writedata),                 //                                 .writedata
		.p1y_s1_chipselect                      (mm_interconnect_0_p1y_s1_chipselect),                //                                 .chipselect
		.p2x_s1_address                         (mm_interconnect_0_p2x_s1_address),                   //                           p2x_s1.address
		.p2x_s1_write                           (mm_interconnect_0_p2x_s1_write),                     //                                 .write
		.p2x_s1_readdata                        (mm_interconnect_0_p2x_s1_readdata),                  //                                 .readdata
		.p2x_s1_writedata                       (mm_interconnect_0_p2x_s1_writedata),                 //                                 .writedata
		.p2x_s1_chipselect                      (mm_interconnect_0_p2x_s1_chipselect),                //                                 .chipselect
		.p2y_s1_address                         (mm_interconnect_0_p2y_s1_address),                   //                           p2y_s1.address
		.p2y_s1_write                           (mm_interconnect_0_p2y_s1_write),                     //                                 .write
		.p2y_s1_readdata                        (mm_interconnect_0_p2y_s1_readdata),                  //                                 .readdata
		.p2y_s1_writedata                       (mm_interconnect_0_p2y_s1_writedata),                 //                                 .writedata
		.p2y_s1_chipselect                      (mm_interconnect_0_p2y_s1_chipselect),                //                                 .chipselect
		.player1_s1_address                     (mm_interconnect_0_player1_s1_address),               //                       player1_s1.address
		.player1_s1_readdata                    (mm_interconnect_0_player1_s1_readdata),              //                                 .readdata
		.player_2_s1_address                    (mm_interconnect_0_player_2_s1_address),              //                      player_2_s1.address
		.player_2_s1_readdata                   (mm_interconnect_0_player_2_s1_readdata),             //                                 .readdata
		.start_s1_address                       (mm_interconnect_0_start_s1_address),                 //                         start_s1.address
		.start_s1_readdata                      (mm_interconnect_0_start_s1_readdata)                 //                                 .readdata
	);

	nios_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
